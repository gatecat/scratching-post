module top(input wire [13:0] A, B, output wire [23:0] X);
	assign X = A*B;
endmodule
